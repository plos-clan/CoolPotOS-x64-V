module storage
