module net
