module hid
