module msc
